`default_nettype none

//分割版

module finv(
	input wire [31:0] x,
        input wire clk,
        input wire rstn,
	output wire [31:0] y);

	wire s;
	wire [7:0] e;
	wire [22:0] m;
	assign {s,e,m} = x;

	wire [23:0] ma;
	assign ma = {1'b1, m};

	function [25:0] INV (
		input [7:0] mh);
	begin
	case (mh)
	8'b00000000: INV = 26'b11111111100000000011111111 ;
        8'b00000001: INV = 26'b11111110100000100011110010 ;
        8'b00000010: INV = 26'b11111101100001100011000010 ;
        8'b00000011: INV = 26'b11111100100011000001010110 ;
        8'b00000100: INV = 26'b11111011100100111110011001 ;
        8'b00000101: INV = 26'b11111010100111011001110100 ;
        8'b00000110: INV = 26'b11111001101010010011010000 ;
        8'b00000111: INV = 26'b11111000101101101010011000 ;
        8'b00001000: INV = 26'b11110111110001011110110110 ;
        8'b00001001: INV = 26'b11110110110101110000010101 ;
        8'b00001010: INV = 26'b11110101111010011110011111 ;
        8'b00001011: INV = 26'b11110100111111101001000010 ;
        8'b00001100: INV = 26'b11110100000101001111100111 ;
        8'b00001101: INV = 26'b11110011001011010001111011 ;
        8'b00001110: INV = 26'b11110010010001101111101011 ;
        8'b00001111: INV = 26'b11110001011000101000100010 ;
        8'b00010000: INV = 26'b11110000011111111100001111 ;
        8'b00010001: INV = 26'b11101111100111101010011110 ;
        8'b00010010: INV = 26'b11101110101111110010111100 ;
        8'b00010011: INV = 26'b11101101111000010101010111 ;
        8'b00010100: INV = 26'b11101101000001010001011110 ;
        8'b00010101: INV = 26'b11101100001010100110111110 ;
        8'b00010110: INV = 26'b11101011010100010101100110 ;
        8'b00010111: INV = 26'b11101010011110011101000101 ;
        8'b00011000: INV = 26'b11101001101000111101001001 ;
        8'b00011001: INV = 26'b11101000110011110101100010 ;
        8'b00011010: INV = 26'b11100111111111000110000000 ;
        8'b00011011: INV = 26'b11100111001010101110010001 ;
        8'b00011100: INV = 26'b11100110010110101110000111 ;
        8'b00011101: INV = 26'b11100101100011000101010001 ;
        8'b00011110: INV = 26'b11100100101111110011011111 ;
        8'b00011111: INV = 26'b11100011111100111000100010 ;
        8'b00100000: INV = 26'b11100011001010010100001011 ;
        8'b00100001: INV = 26'b11100010011000000110001100 ;
        8'b00100010: INV = 26'b11100001100110001110010100 ;
        8'b00100011: INV = 26'b11100000110100101100010110 ;
        8'b00100100: INV = 26'b11100000000011100000000011 ;
        8'b00100101: INV = 26'b11011111010010101001001101 ;
        8'b00100110: INV = 26'b11011110100010000111100110 ;
        8'b00100111: INV = 26'b11011101110001111011000001 ;
        8'b00101000: INV = 26'b11011101000010000011001111 ;
        8'b00101001: INV = 26'b11011100010010100000000011 ;
        8'b00101010: INV = 26'b11011011100011010001010000 ;
        8'b00101011: INV = 26'b11011010110100010110101001 ;
        8'b00101100: INV = 26'b11011010000101110000000001 ;
        8'b00101101: INV = 26'b11011001010111011101001011 ;
        8'b00101110: INV = 26'b11011000101001011101111011 ;
        8'b00101111: INV = 26'b11010111111011110010000101 ;
        8'b00110000: INV = 26'b11010111001110011001011011 ;
        8'b00110001: INV = 26'b11010110100001010011110011 ;
        8'b00110010: INV = 26'b11010101110100100000111111 ;
        8'b00110011: INV = 26'b11010101001000000000110101 ;
        8'b00110100: INV = 26'b11010100011011110011001000 ;
        8'b00110101: INV = 26'b11010011101111110111101110 ;
        8'b00110110: INV = 26'b11010011000100001110011011 ;
        8'b00110111: INV = 26'b11010010011000110111000100 ;
        8'b00111000: INV = 26'b11010001101101110001011101 ;
        8'b00111001: INV = 26'b11010001000010111101011100 ;
        8'b00111010: INV = 26'b11010000011000011010110111 ;
        8'b00111011: INV = 26'b11001111101110001001100010 ;
        8'b00111100: INV = 26'b11001111000100001001010011 ;
        8'b00111101: INV = 26'b11001110011010011010000000 ;
        8'b00111110: INV = 26'b11001101110000111011011110 ;
        8'b00111111: INV = 26'b11001101000111101101100100 ;
        8'b01000000: INV = 26'b11001100011110110000000111 ;
        8'b01000001: INV = 26'b11001011110110000010111111 ;
        8'b01000010: INV = 26'b11001011001101100110000000 ;
        8'b01000011: INV = 26'b11001010100101011001000001 ;
        8'b01000100: INV = 26'b11001001111101011011111010 ;
        8'b01000101: INV = 26'b11001001010101101110100000 ;
        8'b01000110: INV = 26'b11001000101110010000101010 ;
        8'b01000111: INV = 26'b11001000000111000010001111 ;
        8'b01001000: INV = 26'b11000111100000000011000111 ;
        8'b01001001: INV = 26'b11000110111001010011001000 ;
        8'b01001010: INV = 26'b11000110010010110010001001 ;
        8'b01001011: INV = 26'b11000101101100100000000011 ;
        8'b01001100: INV = 26'b11000101000110011100101011 ;
        8'b01001101: INV = 26'b11000100100000100111111010 ;
        8'b01001110: INV = 26'b11000011111011000001101000 ;
        8'b01001111: INV = 26'b11000011010101101001101011 ;
        8'b01010000: INV = 26'b11000010110000011111111100 ;
        8'b01010001: INV = 26'b11000010001011100100010100 ;
        8'b01010010: INV = 26'b11000001100110110110101001 ;
        8'b01010011: INV = 26'b11000001000010010110110011 ;
        8'b01010100: INV = 26'b11000000011110000100101100 ;
        8'b01010101: INV = 26'b10111111111010000000001011 ;
        8'b01010110: INV = 26'b10111111010110001001001001 ;
        8'b01010111: INV = 26'b10111110110010011111011111 ;
        8'b01011000: INV = 26'b10111110001111000011000100 ;
        8'b01011001: INV = 26'b10111101101011110011110001 ;
        8'b01011010: INV = 26'b10111101001000110001100000 ;
        8'b01011011: INV = 26'b10111100100101111100001000 ;
        8'b01011100: INV = 26'b10111100000011010011100011 ;
        8'b01011101: INV = 26'b10111011100000110111101010 ;
        8'b01011110: INV = 26'b10111010111110101000010110 ;
        8'b01011111: INV = 26'b10111010011100100101100000 ;
        8'b01100000: INV = 26'b10111001111010101111000001 ;
        8'b01100001: INV = 26'b10111001011001000100110011 ;
        8'b01100010: INV = 26'b10111000110111100110101110 ;
        8'b01100011: INV = 26'b10111000010110010100101101 ;
        8'b01100100: INV = 26'b10110111110101001110101000 ;
        8'b01100101: INV = 26'b10110111010100010100011010 ;
        8'b01100110: INV = 26'b10110110110011100101111011 ;
        8'b01100111: INV = 26'b10110110010011000011000111 ;
        8'b01101000: INV = 26'b10110101110010101011110110 ;
        8'b01101001: INV = 26'b10110101010010100000000010 ;
        8'b01101010: INV = 26'b10110100110010011111100110 ;
        8'b01101011: INV = 26'b10110100010010101010011011 ;
        8'b01101100: INV = 26'b10110011110011000000011100 ;
        8'b01101101: INV = 26'b10110011010011100001100010 ;
        8'b01101110: INV = 26'b10110010110100001101100111 ;
        8'b01101111: INV = 26'b10110010010101000100100111 ;
        8'b01110000: INV = 26'b10110001110110000110011011 ;
        8'b01110001: INV = 26'b10110001010111010010111101 ;
        8'b01110010: INV = 26'b10110000111000101010001001 ;
        8'b01110011: INV = 26'b10110000011010001011111000 ;
        8'b01110100: INV = 26'b10101111111011111000000110 ;
        8'b01110101: INV = 26'b10101111011101101110101100 ;
        8'b01110110: INV = 26'b10101110111111101111100110 ;
        8'b01110111: INV = 26'b10101110100001111010101101 ;
        8'b01111000: INV = 26'b10101110000100001111111110 ;
        8'b01111001: INV = 26'b10101101100110101111010011 ;
        8'b01111010: INV = 26'b10101101001001011000100110 ;
        8'b01111011: INV = 26'b10101100101100001011110011 ;
        8'b01111100: INV = 26'b10101100001111001000110101 ;
        8'b01111101: INV = 26'b10101011110010001111100110 ;
        8'b01111110: INV = 26'b10101011010101100000000010 ;
        8'b01111111: INV = 26'b10101010111000111010000100 ;
        8'b10000000: INV = 26'b10101010011100011101101000 ;
        8'b10000001: INV = 26'b10101010000000001010101000 ;
        8'b10000010: INV = 26'b10101001100100000000111111 ;
        8'b10000011: INV = 26'b10101001001000000000101010 ;
        8'b10000100: INV = 26'b10101000101100001001100011 ;
        8'b10000101: INV = 26'b10101000010000011011100110 ;
        8'b10000110: INV = 26'b10100111110100110110101111 ;
        8'b10000111: INV = 26'b10100111011001011010111001 ;
        8'b10001000: INV = 26'b10100110111110000111111111 ;
        8'b10001001: INV = 26'b10100110100010111101111101 ;
        8'b10001010: INV = 26'b10100110000111111100110000 ;
        8'b10001011: INV = 26'b10100101101101000100010010 ;
        8'b10001100: INV = 26'b10100101010010010100011111 ;
        8'b10001101: INV = 26'b10100100110111101101010100 ;
        8'b10001110: INV = 26'b10100100011101001110101100 ;
        8'b10001111: INV = 26'b10100100000010111000100011 ;
        8'b10010000: INV = 26'b10100011101000101010110100 ;
        8'b10010001: INV = 26'b10100011001110100101011101 ;
        8'b10010010: INV = 26'b10100010110100101000011000 ;
        8'b10010011: INV = 26'b10100010011010110011100011 ;
        8'b10010100: INV = 26'b10100010000001000110111000 ;
        8'b10010101: INV = 26'b10100001100111100010010100 ;
        8'b10010110: INV = 26'b10100001001110000101110100 ;
        8'b10010111: INV = 26'b10100000110100110001010100 ;
        8'b10011000: INV = 26'b10100000011011100100101111 ;
        8'b10011001: INV = 26'b10100000000010100000000010 ;
        8'b10011010: INV = 26'b10011111101001100011001010 ;
        8'b10011011: INV = 26'b10011111010000101110000010 ;
        8'b10011100: INV = 26'b10011110111000000000100111 ;
        8'b10011101: INV = 26'b10011110011111011010110110 ;
        8'b10011110: INV = 26'b10011110000110111100101011 ;
        8'b10011111: INV = 26'b10011101101110100110000010 ;
        8'b10100000: INV = 26'b10011101010110010110111001 ;
        8'b10100001: INV = 26'b10011100111110001111001011 ;
        8'b10100010: INV = 26'b10011100100110001110110101 ;
        8'b10100011: INV = 26'b10011100001110010101110100 ;
        8'b10100100: INV = 26'b10011011110110100100000100 ;
        8'b10100101: INV = 26'b10011011011110111001100010 ;
        8'b10100110: INV = 26'b10011011000111010110001100 ;
        8'b10100111: INV = 26'b10011010101111111001111101 ;
        8'b10101000: INV = 26'b10011010011000100100110010 ;
        8'b10101001: INV = 26'b10011010000001010110101000 ;
        8'b10101010: INV = 26'b10011001101010001111011101 ;
        8'b10101011: INV = 26'b10011001010011001111001100 ;
        8'b10101100: INV = 26'b10011000111100010101110011 ;
        8'b10101101: INV = 26'b10011000100101100011001111 ;
        8'b10101110: INV = 26'b10011000001110110111011100 ;
        8'b10101111: INV = 26'b10010111111000010010011001 ;
        8'b10110000: INV = 26'b10010111100001110100000000 ;
        8'b10110001: INV = 26'b10010111001011011100010001 ;
        8'b10110010: INV = 26'b10010110110101001011000111 ;
        8'b10110011: INV = 26'b10010110011111000000100000 ;
        8'b10110100: INV = 26'b10010110001000111100011010 ;
        8'b10110101: INV = 26'b10010101110010111110110000 ;
        8'b10110110: INV = 26'b10010101011101000111100001 ;
        8'b10110111: INV = 26'b10010101000111010110101001 ;
        8'b10111000: INV = 26'b10010100110001101100000110 ;
        8'b10111001: INV = 26'b10010100011100000111110100 ;
        8'b10111010: INV = 26'b10010100000110101001110011 ;
        8'b10111011: INV = 26'b10010011110001010001111101 ;
        8'b10111100: INV = 26'b10010011011100000000010010 ;
        8'b10111101: INV = 26'b10010011000110110100101110 ;
        8'b10111110: INV = 26'b10010010110001101111001110 ;
        8'b10111111: INV = 26'b10010010011100101111110001 ;
        8'b11000000: INV = 26'b10010010000111110110010010 ;
        8'b11000001: INV = 26'b10010001110011000010110001 ;
        8'b11000010: INV = 26'b10010001011110010101001010 ;
        8'b11000011: INV = 26'b10010001001001101101011011 ;
        8'b11000100: INV = 26'b10010000110101001011100001 ;
        8'b11000101: INV = 26'b10010000100000101111011010 ;
        8'b11000110: INV = 26'b10010000001100011001000100 ;
        8'b11000111: INV = 26'b10001111111000001000011011 ;
        8'b11001000: INV = 26'b10001111100011111101011110 ;
        8'b11001001: INV = 26'b10001111001111111000001010 ;
        8'b11001010: INV = 26'b10001110111011111000011101 ;
        8'b11001011: INV = 26'b10001110100111111110010101 ;
        8'b11001100: INV = 26'b10001110010100001001101110 ;
        8'b11001101: INV = 26'b10001110000000011010101000 ;
        8'b11001110: INV = 26'b10001101101100110000111111 ;
        8'b11001111: INV = 26'b10001101011001001100110001 ;
        8'b11010000: INV = 26'b10001101000101101101111100 ;
        8'b11010001: INV = 26'b10001100110010010100011111 ;
        8'b11010010: INV = 26'b10001100011111000000010101 ;
        8'b11010011: INV = 26'b10001100001011110001011111 ;
        8'b11010100: INV = 26'b10001011111000100111111000 ;
        8'b11010101: INV = 26'b10001011100101100011100000 ;
        8'b11010110: INV = 26'b10001011010010100100010100 ;
        8'b11010111: INV = 26'b10001010111111101010010010 ;
        8'b11011000: INV = 26'b10001010101100110101010111 ;
        8'b11011001: INV = 26'b10001010011010000101100010 ;
        8'b11011010: INV = 26'b10001010000111011010110001 ;
        8'b11011011: INV = 26'b10001001110100110101000001 ;
        8'b11011100: INV = 26'b10001001100010010100010001 ;
        8'b11011101: INV = 26'b10001001001111111000011111 ;
        8'b11011110: INV = 26'b10001000111101100001101000 ;
        8'b11011111: INV = 26'b10001000101011001111101011 ;
        8'b11100000: INV = 26'b10001000011001000010100110 ;
        8'b11100001: INV = 26'b10001000000110111010010110 ;
        8'b11100010: INV = 26'b10000111110100110110111010 ;
        8'b11100011: INV = 26'b10000111100010111000010000 ;
        8'b11100100: INV = 26'b10000111010000111110010110 ;
        8'b11100101: INV = 26'b10000110111111001001001010 ;
        8'b11100110: INV = 26'b10000110101101011000101010 ;
        8'b11100111: INV = 26'b10000110011011101100110101 ;
        8'b11101000: INV = 26'b10000110001010000101101000 ;
        8'b11101001: INV = 26'b10000101111000100011000010 ;
        8'b11101010: INV = 26'b10000101100111000101000001 ;
        8'b11101011: INV = 26'b10000101010101101011100011 ;
        8'b11101100: INV = 26'b10000101000100010110100111 ;
        8'b11101101: INV = 26'b10000100110011000110001010 ;
        8'b11101110: INV = 26'b10000100100001111010001011 ;
        8'b11101111: INV = 26'b10000100010000110010101000 ;
        8'b11110000: INV = 26'b10000011111111101111100000 ;
        8'b11110001: INV = 26'b10000011101110110000110000 ;
        8'b11110010: INV = 26'b10000011011101110110010111 ;
        8'b11110011: INV = 26'b10000011001101000000010100 ;
        8'b11110100: INV = 26'b10000010111100001110100100 ;
        8'b11110101: INV = 26'b10000010101011100001000111 ;
        8'b11110110: INV = 26'b10000010011010110111111010 ;
        8'b11110111: INV = 26'b10000010001010010010111100 ;
        8'b11111000: INV = 26'b10000001111001110010001011 ;
        8'b11111001: INV = 26'b10000001101001010101100101 ;
        8'b11111010: INV = 26'b10000001011000111101001010 ;
        8'b11111011: INV = 26'b10000001001000101000110110 ;
        8'b11111100: INV = 26'b10000000111000011000101010 ;
        8'b11111101: INV = 26'b10000000101000001100100011 ;
        8'b11111110: INV = 26'b10000000011000000100100000 ;
        8'b11111111: INV = 26'b10000000001000000000100000;
	default : INV = 26'bx;
	endcase
	end
	endfunction

	wire [25:0] init;
	assign init = INV(ma[22:15]);

	wire [74:0] k1;
 	assign k1 = {51'b0, ma} * {49'b0, init} * {49'b0, init};

        logic [23:0] ma1;
        logic [25:0] init1;
        logic [74:0] k11;
        logic s1;
        logic [7:0] e1;

        always @(posedge clk) begin
                ma1 <= ma;
                init1 <= init;
                k11 <= k1;
                s1 <= s;
                e1 <= e;
        end

 	wire [75:0] c1;
 	assign c1 = {init1, 50'b0} - {1'b0, k11};

 	wire [25:0] x1;
 	assign x1 = (c1[48] && (|c1[47:0] || c1[49]))? {c1[74:49]} + 26'b1
 						: {c1[74:49]};

        logic [23:0] ma2;
        logic [25:0] x11;
        logic s2;
        logic [7:0] e2;

        always @(posedge clk) begin
                ma2 <= ma1;
                x11 <= x1;
                s2 <= s1;
                e2 <= e1;
        end

 	wire [74:0] k2;
 	assign k2 = {51'b0, ma2} * {49'b0, x11} * {49'b0, x11};

 	wire [75:0] c2;
 	assign c2 = {x11, 50'b0} - {1'b0, k2};

 	wire [25:0] x2;
 	assign x2 = (c2[48] && (|c2[47:0] || c2[49]))? {c2[74:49]} + 26'b1
 							: {c2[74:49]};

 	wire [7:0] ey;
 	wire [22:0] my;

 	assign my = (e2 == 8'd254)? ((x2[3])? {1'b0, x2[25:4]} + 23'b1
 					: {1'b0, x2[25:4]}) 
                                        :(e2 == 8'd253)? ((x2[2])? x2[25:3] + 23'b1 : x2[25:3]) 
                                        :(x2[1])? x2[24:2] + 23'b1 : x2[24:2];

 	assign ey = (e2 == 8'd254)? ~e2 - 1: ~e2 - 2;

 	assign y = (my == 23'b0) ? {s2,ey + 8'b1, my} : {s2,ey,my};

 endmodule

 `default_nettype wire