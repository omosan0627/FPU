`default_nettype none

module fsqrt(
  input wire [31:0] x,
  output wire [31:0] y);

  wire s;
  wire [7:0] e;
  wire [22:0] m;

  assign {s,e,m} = x;

  wire [24:0] ma;
  assign ma =  (|e && ~e[0:0]) ? {2'b1,m} :
                (|e && e[0:0]) ? {1'b1,m,1'b0} :
                (m[22]) ? {1'b0,m,1'b0} :
                (m[21] || m[20]) ? {m[21:0],3'b0} :
                (m[19] || m[18]) ? {m[19:0],5'b0} : 
                (m[17] || m[16]) ? {m[17:0],7'b0} : 
                (m[15] || m[14]) ? {m[15:0],9'b0} : 
                (m[13] || m[12]) ? {m[13:0],11'b0} : 
                (m[11] || m[10]) ? {m[11:0],13'b0} : 
                (m[9] || m[8]) ? {m[9:0],15'b0} : 
                (m[7] || m[6]) ? {m[7:0],17'b0} : 
                (m[5] || m[4]) ? {m[5:0],19'b0} : 
                (m[3] || m[2]) ? {m[3:0],21'b0} : {m[1:0],23'b0};

  wire [7:0] ea;
  assign ea = (|e) ? {1'b0,e[7:1]} + 64 :
               (m[22]) ? 8'd64 :
               (m[21] || m[20]) ? 63 :
               (m[19] || m[18]) ? 62 : 
               (m[17] || m[16]) ? 61 : 
               (m[15] || m[14]) ? 60 : 
               (m[13] || m[12]) ? 59 : 
               (m[11] || m[10]) ? 58 : 
               (m[9] || m[8]) ? 57 : 
               (m[7] || m[6]) ? 56 : 
               (m[5] || m[4]) ? 55 : 
               (m[3] || m[2]) ? 54 : 53;

  wire [27:0] init;
  assign init = {2'b1, 26'b0};

  wire [27:0] y1;
  wire [106:0] p1;
  assign p1 = ({27'b0,2'b11,78'b0} - ({80'b0,ma,2'b0} * {79'b0,init} * {79'b0,init})) * {79'b0,init};
  assign y1 = (p1[78] && (|p1[77:0] || p1[79])) ? p1[106:79] + 28'b1 : p1[106:79];

  wire [27:0] y2;
  wire [106:0] p2;
  assign p2 = ({27'b0,2'b11,78'b0} - ({80'b0,ma,2'b0} * {79'b0,y1} * {79'b0,y1})) * {79'b0,y1};
  assign y2 = (p2[78] && (|p2[77:0] || p2[79])) ? p2[106:79] + 28'b1 : p2[106:79];

  wire [27:0] y3;
  wire [106:0] p3;
  assign p3 = ({27'b0,2'b11,78'b0} - ({80'b0,ma,2'b0} * {79'b0,y2} * {79'b0,y2})) * {79'b0,y2};
  assign y3 = (p3[78] && (|p3[77:0] || p3[79])) ? p3[106:79] + 28'b1 : p3[106:79];

  wire [27:0] y4;
  wire [106:0] p4;
  assign p4 = ({27'b0,2'b11,78'b0} - ({80'b0,ma,2'b0} * {79'b0,y3} * {79'b0,y3})) * {79'b0,y3};
  assign y4 = (p4[78] && (|p4[77:0] || p4[79])) ? p4[106:79] + 28'b1 : p4[106:79];

  wire [27:0] y5;
  wire [106:0] p5;
  assign p5 = ({27'b0,2'b11,78'b0} - ({80'b0,ma,2'b0} * {79'b0,y4} * {79'b0,y4})) * {79'b0,y4};
  assign y5 = (p5[78] && (|p5[77:0] || p5[79])) ? p5[106:79] + 28'b1 : p5[106:79];

  wire [24:0] mye;
  assign mye = (y5[27]) ? ((y5[3]) ? {1'b0, y5[27:4]} + 25'b1 : {1'b0, y5[27:4]}) :
                (y5[26]) ? ((y5[2]) ? {1'b0, y5[26:3]} + 25'b1 : {1'b0, y5[26:3]}) :
                (y5[25]) ? ((y5[1]) ? {1'b0, y5[25:2]} + 25'b1 : {1'b0, y5[25:2]}) :
                (y5[0]) ? {1'b0, y5[24:1]} + 25'b0 : {1'b0, y5[24:1]};

  wire [22:0] my;
  assign my = (mye[24]) ? 23'b0 : mye[22:0];

  wire [7:0] eye;
  assign eye = (y5[27]) ? 255 - ea :
                (y5[26]) ? 254 - ea :
                (y5[25]) ? 253 - ea : 252 - ea;

  wire [7:0] ey;
  assign ey = (mye[24]) ? eye + 8'b1 : eye;

  wire [31:0] y_mul;
  wire ovf_mul;

  fmul u1(x, {s, ey, my}, y_mul, ovf_mul);

  wire nzm;
  assign nzm = |m;

  assign y =  (e == 8'd255 && nzm) ? {s,8'd255,1'b1,m[21:0]} : 
              (s == 1'b0 && e == 8'd255 && ~nzm) ? {1'b0,8'd255,23'b0} :
              (~|x) ? {1'b0,8'b0,23'b0} : 
              (s == 1'b1 && ~|x[30:0]) ? {1'b1,8'b0,23'b0} : 
              (s == 1'b1) ? {1'b1,8'd255,1'b1,22'b0} : y_mul;
endmodule

`default_nettype wire